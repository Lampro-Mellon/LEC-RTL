#(parameter
	 AWIDTH = 7,
	 TAG = 1'h1,
	 BHT_ADDR_HI =  4'h9 ,
	 BHT_ADDR_LO =  2'h2 ,
	 BHT_ARRAY_DEPTH =  11'h100 ,
	 BHT_GHR_HASH_1 =  1'h0 ,
	 BHT_GHR_SIZE =  4'h8 ,
	 BHT_SIZE =  12'h200 ,
	 BTB_ADDR_HI =  5'h09 ,
	 BTB_ADDR_LO =  2'h2 ,
	 BTB_ARRAY_DEPTH =  9'h100 ,
	 BTB_BTAG_FOLD =  1'h0 ,
	 BTB_BTAG_SIZE =  4'h5 ,
	 BTB_FOLD2_INDEX_HASH =  1'h0 ,
	 BTB_INDEX1_HI =  5'h09 ,
	 BTB_INDEX1_LO =  5'h02 ,
	 BTB_INDEX2_HI =  5'h11 ,
	 BTB_INDEX2_LO =  5'h0A ,
	 BTB_INDEX3_HI =  5'h19 ,
	 BTB_INDEX3_LO =  5'h12 ,
	 BTB_SIZE =  10'h200 ,
	 BUILD_AHB_LITE =  1'h0 ,
	 BUILD_AXI4 =  1'h1 ,
	 BUILD_AXI_NATIVE =  1'h1 ,
	 BUS_PRTY_DEFAULT =  2'h3 ,
	 DATA_ACCESS_ADDR0 =  32'h00000000 ,
	 DATA_ACCESS_ADDR1 =  32'hC0000000 ,
	 DATA_ACCESS_ADDR2 =  32'hA0000000 ,
	 DATA_ACCESS_ADDR3 =  32'h80000000 ,
	 DATA_ACCESS_ADDR4 =  32'h00000000 ,
	 DATA_ACCESS_ADDR5 =  32'h00000000 ,
	 DATA_ACCESS_ADDR6 =  32'h00000000 ,
	 DATA_ACCESS_ADDR7 =  32'h00000000 ,
	 DATA_ACCESS_ENABLE0 =  1'h1 ,
	 DATA_ACCESS_ENABLE1 =  1'h1 ,
	 DATA_ACCESS_ENABLE2 =  1'h1 ,
	 DATA_ACCESS_ENABLE3 =  1'h1 ,
	 DATA_ACCESS_ENABLE4 =  1'h0 ,
	 DATA_ACCESS_ENABLE5 =  1'h0 ,
	 DATA_ACCESS_ENABLE6 =  1'h0 ,
	 DATA_ACCESS_ENABLE7 =  1'h0 ,
	 DATA_ACCESS_MASK0 =  32'h7FFFFFFF ,
	 DATA_ACCESS_MASK1 =  32'h3FFFFFFF ,
	 DATA_ACCESS_MASK2 =  32'h1FFFFFFF ,
	 DATA_ACCESS_MASK3 =  32'h0FFFFFFF ,
	 DATA_ACCESS_MASK4 =  32'hFFFFFFFF ,
	 DATA_ACCESS_MASK5 =  32'hFFFFFFFF ,
	 DATA_ACCESS_MASK6 =  32'hFFFFFFFF ,
	 DATA_ACCESS_MASK7 =  32'hFFFFFFFF ,
	 DCCM_BANK_BITS =  3'h2 ,
	 DCCM_BITS =  5'h11 ,
	 DCCM_BYTE_WIDTH =  3'h4 ,
	 DCCM_DATA_WIDTH =  6'h20 ,
	 DCCM_ECC_WIDTH =  3'h7 ,
	 DCCM_ENABLE =  1'h1 ,
	 DCCM_FDATA_WIDTH =  6'h27 ,
	// DCCM_INDEX_BITS =  4'hC ,
	 DCCM_NUM_BANKS =  5'h04 ,
	 DCCM_REGION =  4'hF ,
	 DCCM_SADR =  32'hF0040000 ,
	 DCCM_SIZE =  10'h080 ,
	 DCCM_WIDTH_BITS =  2'h2 ,
	 DMA_BUF_DEPTH =  3'h5 ,
	 DMA_BUS_ID =  1'h1 ,
	 DMA_BUS_PRTY =  2'h2 ,
	 DMA_BUS_TAG =  4'h1 ,
	 FAST_INTERRUPT_REDIRECT =  1'h1 ,
	 ICACHE_2BANKS =  1'h1 ,
	 ICACHE_BANK_BITS =  3'h1 ,
	 ICACHE_BANK_HI =  3'h3 ,
	 ICACHE_BANK_LO =  2'h3 ,
	 ICACHE_BANK_WIDTH =  4'h8 ,
	 ICACHE_BANKS_WAY =  3'h2 ,
	 ICACHE_BEAT_ADDR_HI =  4'h5 ,
	 ICACHE_BEAT_BITS =  4'h3 ,
	 ICACHE_DATA_DEPTH =  14'h0200 ,
	 ICACHE_DATA_INDEX_LO =  3'h4 ,
	 ICACHE_DATA_WIDTH =  7'h40 ,
	 ICACHE_ECC =  1'h1 ,
	 ICACHE_ENABLE =  1'h1 ,
	 ICACHE_FDATA_WIDTH =  7'h47 ,
	 ICACHE_INDEX_HI =  5'h0C ,
	 ICACHE_LN_SZ =  7'h40 ,
	 ICACHE_NUM_BEATS =  4'h8 ,
	 ICACHE_NUM_WAYS =  3'h2 ,
	 ICACHE_ONLY =  1'h0 ,
	 ICACHE_SCND_LAST =  4'h6 ,
	 ICACHE_SIZE =  9'h010 ,
	 ICACHE_STATUS_BITS =  3'h1 ,
	 ICACHE_TAG_DEPTH =  13'h0080 ,
	 ICACHE_TAG_INDEX_LO =  3'h6 ,
	 ICACHE_TAG_LO =  5'h0D ,
	 ICACHE_WAYPACK =  1'h0 ,
	 ICCM_BANK_BITS =  3'h2 ,
	 ICCM_BANK_HI =  5'h03 ,
	 ICCM_BANK_INDEX_LO =  5'h04 ,
	 ICCM_BITS =  5'h10 ,
	 ICCM_ENABLE =  1'h1 ,
	 ICCM_ICACHE =  1'h1 ,
	 ICCM_INDEX_BITS =  4'hC ,
	 ICCM_NUM_BANKS =  5'h04 ,
	 ICCM_ONLY =  1'h0 ,
	 ICCM_REGION =  4'hE ,
	 ICCM_SADR =  32'hEE000000 ,
	 ICCM_SIZE =  10'h040 ,
	 IFU_BUS_ID =  1'h1 ,
	 IFU_BUS_PRTY =  2'h2 ,
	 IFU_BUS_TAG =  4'h3 ,
	 INST_ACCESS_ADDR0 =  32'h00000000 ,
	 INST_ACCESS_ADDR1 =  32'hC0000000 ,
	 INST_ACCESS_ADDR2 =  32'hA0000000 ,
	 INST_ACCESS_ADDR3 =  32'h80000000 ,
	 INST_ACCESS_ADDR4 =  32'h00000000 ,
	 INST_ACCESS_ADDR5 =  32'h00000000 ,
	 INST_ACCESS_ADDR6 =  32'h00000000 ,
	 INST_ACCESS_ADDR7 =  32'h00000000 ,
	 INST_ACCESS_ENABLE0 =  1'h1 ,
	 INST_ACCESS_ENABLE1 =  1'h1 ,
	 INST_ACCESS_ENABLE2 =  1'h1 ,
	 INST_ACCESS_ENABLE3 =  1'h1 ,
	 INST_ACCESS_ENABLE4 =  1'h0 ,
	 INST_ACCESS_ENABLE5 =  1'h0 ,
	 INST_ACCESS_ENABLE6 =  1'h0 ,
	 INST_ACCESS_ENABLE7 =  1'h0 ,
	 INST_ACCESS_MASK0 =  32'h7FFFFFFF ,
	 INST_ACCESS_MASK1 =  32'h3FFFFFFF ,
	 INST_ACCESS_MASK2 =  32'h1FFFFFFF ,
	 INST_ACCESS_MASK3 =  32'h0FFFFFFF ,
	 INST_ACCESS_MASK4 =  32'hFFFFFFFF ,
	 INST_ACCESS_MASK5 =  32'hFFFFFFFF ,
	 INST_ACCESS_MASK6 =  32'hFFFFFFFF ,
	 INST_ACCESS_MASK7 =  32'hFFFFFFFF ,
	 LOAD_TO_USE_PLUS1 =  1'h0 ,
	 LSU2DMA =  1'h0 ,
	 LSU_BUS_ID =  1'h1 ,
	 LSU_BUS_PRTY =  2'h2 ,
	 LSU_BUS_TAG =  4'h3 ,
	 LSU_NUM_NBLOAD =  5'h04 ,
	 LSU_NUM_NBLOAD_WIDTH =  3'h2 ,
	 LSU_SB_BITS =  5'h11 ,
	 LSU_STBUF_DEPTH =  4'h4 ,
	 NO_ICCM_NO_ICACHE =  1'h0 ,
	 PIC_2CYCLE =  1'h0 ,
	 PIC_BASE_ADDR =  32'hF00C0000 ,
	 PIC_BITS =  5'h0F ,
	 PIC_INT_WORDS =  4'h1 ,
	 PIC_REGION =  4'hF ,
	 PIC_SIZE =  9'h020 ,
	 PIC_TOTAL_INT =  8'h1F ,
	 PIC_TOTAL_INT_PLUS1 =  9'h020 ,
	 RET_STACK_SIZE =  4'h8 ,
	 SB_BUS_ID =  1'h1 ,
	 SB_BUS_PRTY =  2'h2 ,
	 SB_BUS_TAG =  4'h1 ,
	 TIMER_LEGAL_EN =  1'h1
)
